library verilog;
use verilog.vl_types.all;
entity Proj_rev2_vlg_vec_tst is
end Proj_rev2_vlg_vec_tst;
